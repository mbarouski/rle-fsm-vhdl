-------------------------------------------------------------------------------
--
-- Title       : GPR_UNIT_X
-- Design      : fsm_rle
-- Author      : maxim
-- Company     : none
--
-------------------------------------------------------------------------------
--
-- File        : GPR_UNIT_X.vhd
-- Generated   : Sat Nov 30 13:57:17 2019
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {GPR_UNIT_X} architecture {GPR_UNIT_X}}

library IEEE;
use IEEE.STD_LOGIC_1164.all; 
use FSM_RLE.all;

entity GPR_UNIT_X is 
	port(
		GPR_IN : in GPR_UNIT_OUTPUTS;
		GPR_OUT : out GPR_UNIT_INPUTS
		);
end GPR_UNIT_X;

--}} End of automatically maintained section

architecture GPR_UNIT_X of GPR_UNIT_X is
begin

	 -- enter your statements here --

end GPR_UNIT_X;
