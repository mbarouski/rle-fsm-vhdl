-------------------------------------------------------------------------------
--
-- Title       : RAM_UNIT_X
-- Design      : fsm_rle
-- Author      : maxim
-- Company     : none
--
-------------------------------------------------------------------------------
--
-- File        : RAM_UNIT_X.vhd
-- Generated   : Sat Nov 30 13:00:07 2019
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

library IEEE;				 			
use IEEE.STD_LOGIC_1164.all;
use FSM_RLE.all;

entity RAM_UNIT_X is
	port(
		RAM_IN : in RAM_UNIT_OUTPUTS;
		RAM_OUT : out RAM_UNIT_INPUTS
		);
end RAM_UNIT_X;							

architecture RAM_UNIT_X of RAM_UNIT_X is 
	
	--component RAM_UNIT is
--		port(
--			CLK : in STD_LOGIC;
--			RST : in STD_LOGIC;
--			TOS : in NIBBLE;
--			TOS_1 : in BYTE;
--			IR : in NIBBLE;
--			ADR_SEL : in STD_LOGIC;
--			ADR_EN : in STD_LOGIC;
--			DATA_EN : in STD_LOGIC;
--			W_EN : in STD_LOGIC;
--			R_EN : in STD_LOGIC;
--			RAM_DATA : out BYTE
--			);
--	end component;
	
begin
	
	-- enter your statements here --
	
end RAM_UNIT_X;
